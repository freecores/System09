--==========================================================================--
--                                                                          --
-- Synthesizable SYS09BUG Monitor Program for XESS XSA-3S1000 & XuLA boards --
--                                                                          --
--==========================================================================--
--
--  File name      : sys09bug_xes_rom4k_b16.vhd
--
--  Entity name    : mon_rom
--
--  Purpose        : Implements a 4KByte Sys09bug monitor ROM for System09
--                   as implemented on the XESS XSA-3S1000 & XuLA FPGA boards
--
--  Dependencies   : ieee.std_logic_1164
--                   ieee.std_logic_arith
--
--  Uses           : RAMB16_S9 (Xilinx 16KBit Block RAM)
--
--  Author         : John E. Kent
--
--  Email          : dilbert57@opencores.org      
--
--  Web            : http://opencores.org/project,system09
--
--  Description    : Sys09bug monitor ROM for the XESS XSA-3S1000 and XuLA FPGA Boards
--                   Resides at $F000-$FFFF
--                   The lower 2KB ($F000-$F7FF) is read/writeable
--                   The upper 2KB ($F800-$FFFF) is read only
--                   Assumes I/O   at $E000-$EFFF
--                   Control ACIA  at $E000-$E001
--                   PS/2 keyboard at $E020-$E021
--                   VDU8          at $E030-$E034
--                   IDE interface at $E100-$E13F
--                   Assumes RAM   at $DFC0-$DFFF
--
--  Copyright (C) 2011 John Kent
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--===========================================================================--
--                                                                           --
--                              Revision  History                            --
--                                                                           --
--===========================================================================--
--
-- Version Date        Author     Changes
--
-- 1.0     2006-11-21  John Kent  Initial release
-- 1.1     2006-12-22  John Kent  made into 4K ROM/RAM.
-- 1.2     2011-06-04  John Kent  Updated header and description and added GPL
--                                Made lower 2KB ($F000-$F7FF) read/writeable
--                                Made upper 2KB ($F800-$FFFF) read only
-- 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
library unisim;
	use unisim.vcomponents.all;

entity mon_rom is
    Port (
       clk      : in  std_logic;
		 rst      : in  std_logic;
		 cs       : in  std_logic;
		 rw       : in  std_logic;
       addr     : in  std_logic_vector (11 downto 0);
       data_in  : in  std_logic_vector (7 downto 0);
       data_out : out std_logic_vector (7 downto 0)
    );
end mon_rom;

architecture rtl of mon_rom is

  signal we        : std_logic;
  signal cs0       : std_logic;
  signal cs1       : std_logic;
  signal dp0       : std_logic;
  signal dp1       : std_logic;
  signal data_out0 : std_logic_vector(7 downto 0);
  signal data_out1 : std_logic_vector(7 downto 0);


begin

  --
  -- lower block is writeable
  --
  ROM0 : RAMB16_S9
    generic map ( 
    INIT_00 => x"8C02300D2780E12CF08E20C0022F60C10AF89FAD2086891F7F8406F89FAD02F0",
    INIT_01 => x"CD8E040D0A3F2054414857B7F258E1F0463EF042946E24021635F08EF52635F0",
    INIT_02 => x"B6B035EE261F30F6263F310A254700E0B6E2048E10E8038E30343B341F4AAF00",
    INIT_03 => x"0235ED261F30F5263F310C25474700E0B6E2048E10E8038E02343034B03501E0",
    INIT_04 => x"2E2E2E6B7369642045444920676E6974616D726F460D0AB03501E0B70235B035",
    INIT_05 => x"6E20657669726420454449040D0A043F207265626D754E2065766972440D0A20",
    INIT_06 => x"6574656C706D6F432074616D726F460D0A04202164657461636F6C6C6120746F",
    INIT_07 => x"3080ED0022103381F3002510308172FF17FB2459FF174EF2BD89F08EB8F4BD04",
    INIT_08 => x"00028E0201B7018601017FFB265A80A75F4F00028E35F5BDFD008E0001F7891F",
    INIT_09 => x"B602017C10F5BD0201F60101B601A70186846C042600814C0201B684A70101B6",
    INIT_0a => x"8EECF4BDFFC63F8600028EC82640810101B601017C0201B70186D72600810201",
    INIT_0b => x"FFC64F016F846F00028EECF4BDFFC64F00028E10F5BDFFC63F86016F846F0002",
    INIT_0c => x"CC1288ED444DCC1088ED4152CC016F846F00028EECF4BD03C64F00028E10F5BD",
    INIT_0d => x"88ED1F88EDFFC63F861D88ED0101CC1B88ED0100CC1688ED204BCC1488ED5349",
    INIT_0e => x"4F00F78E10F5BD03C64F2588A707862488A707862388A701862188EDC13ECC26",
    INIT_0f => x"E0B7118600E0B7038639018500E0B64EF27ECFF08E2503170201F70101B701C6",
    INIT_10 => x"1C01E0B6E620DD8D0A2778850826018500E0B60A017F09017F0801B710863900",
    INIT_11 => x"78850826028500E0B6023439021A4FDC2608017AE12609017AE6260A017A39FD",
    INIT_12 => x"4449206D65646F6D580A0D39F826048180A6E78D3901E0B70235F120B38DF527",
    INIT_13 => x"046574656C706D6F432064616F6C70550A0D0464616F6C7055206B7369442045",
    INIT_14 => x"043A207265626D754E2065766972440A0D04726F7272452064616F6C70550A0D",
    INIT_15 => x"8FF28E91FF1755F28E04294E2F5928203F206572755320756F59206572410A0D",
    INIT_16 => x"178FF28E0001B730802801221033812E01251030816AFF17FB293CFF178BFF17",
    INIT_17 => x"FF0027104E815F843DFF17FB290FFF175EFF17A0F28E4BFF17308B0001B66CFF",
    INIT_18 => x"00170201F70101B701C64F00028E0401B701860601FF28F4CEB10117B3265981",
    INIT_19 => x"028E710117D501170201F60101B600028ED6002510E00017870117E0002510EA",
    INIT_1a => x"8EA6002510B00017570117B0002510BA00170201F70101B75C0201F60101B600",
    INIT_1b => x"00170201F70101B75C0201F60101B600028E410117A501170201F60101B60002",
    INIT_1c => x"0C01F75C2788E60B01B74C2688A600028E76002510800017270117800025108A",
    INIT_1d => x"104C00170201F70101B700028E5C0201F60101B60301176701170201F60101B6",
    INIT_1e => x"F60101B6D300173701170201F60101B600028E38002510420017E90017420025",
    INIT_1f => x"8E1101170201F70101B701C64F00F78EC3260B01B14C01C6CB260C01F15C0201",
    INIT_20 => x"ADF12028F4CE1BFE1715860A28EFFD170601FE403443FE1680F28E4EF27E6EF2",
    INIT_21 => x"188139051AFAFD1706860826048139FA1C48F4CE06260181C0350601FFED26C4",
    INIT_22 => x"B14339FA1C28F4CEDDFD17158639FA1C5EF4CE06260401B139FA1C39051A0326",
    INIT_23 => x"2605017A02350301B70301BB023439FA1C72F4CE0501B7808603017FEF260401",
    INIT_24 => x"80C45A101F043439041AFE1C28F4CE04017C0B260301B139FA1C80A789F4CE03",
    INIT_25 => x"00CC1EE1FD0600CC82357FFD170686023439FA1C28F4CE8CFD1715860435011F",
    INIT_26 => x"01F608E1FDE4E606E1FD5A4F023401C64F668DDB02160CE1FDE000CC1EE1FD02",
    INIT_27 => x"B7021700018E102034B102170EE1FD2000CCE48D82355F04E1FD01C60AE1FD00",
    INIT_28 => x"018E1020348D02170EE1FD3000CCC08D395F9A02172035F4263F3180E700E1FC",
    INIT_29 => x"5F0001B74F0123038103A6395F7502172035F4263F3100E1FD80E69202174F00",
    INIT_2a => x"000000000000000000000000000000000000000000000000000000395F03A639",
    INIT_2b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"270281358D00C48E1000C3FDF18CECFFC0CE1000000000C00000000000000B20",
    INIT_39 => x"5D891F158DD08CA71A8DD48CA71F8DEA20DA8CA7268DDE8CA72B8DF626168110",
    INIT_3a => x"8D0B2784EC00C38E0F2600C48C10C920F5265A80A71435098D1434C58CAED927",
    INIT_3b => x"C60AE1FD908CE608E1FDE4E606E1FD5A4F02349B9C6E39A0A604C38E109D2626",
    INIT_3c => x"3F3180E700E1FC1E8D00018E102034178D0EE1FD2000CCE48D82355F04E1FD01",
    INIT_3d => x"0039F92708C50EE1FC39F22740C50EE1FCF92680C50EE1FC395F028D2035F526",
    INIT_3e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3f => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out0,
	  dop(0) => dp0,
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp0,
	  en   => cs0,
	  ssr  => rst,
	  we   => we
	);

  --
  -- upper block is not writeable
  --
  ROM1 : RAMB16_S9
    generic map ( 
    INIT_00 => x"A780A610C6C0DF8E1074FE8E2EFA1AFB1EFB8FFBCEFCB9FC9BFCA1FC61F814F8",
    INIT_01 => x"17431FE4A7D0866AAFDD8C30FB265AE26F0CC65B0117E0DFBF00E08EF9265AA0",
    INIT_02 => x"0317A3FE8E0C0417F62A5A19048B0327856D0DC64FD0DF8E47031784FE8E9F04",
    INIT_03 => x"17408B981F5304175E86092C2081891FF1270D817F84370417B30217AAFE8E2E",
    INIT_04 => x"20F00217ACFE8EF52674FE8C02300F2780E13BFE8E20C0022F60C14704174C04",
    INIT_05 => x"17A4A60F0417A50317211F650217B2FE8E121F2D296B03173B341FBC2094ADC0",
    INIT_06 => x"27A4A1A4A7390F260D8117275E81DD271881E127088111285E0317070417A503",
    INIT_07 => x"0B031705201F30C0DF8E321FA20217BE203F31C2202131E503173F86E8031708",
    INIT_08 => x"279A03170527E4AC011FF0C4201F0634F0C41000C3101F390124E1AC20340629",
    INIT_09 => x"265A8E03172C031780A610C69603172E0317E4AEEE0117B2FE8E103439623203",
    INIT_0a => x"29B70217BC20EE265A7703172E8602237E810425208180A610C6E1AE860317F5",
    INIT_0b => x"3984A73F86A4AFA0A709273F8184A60F271035558DFFFF8E10341A24C0DF8C1E",
    INIT_0c => x"4AAF0427268D1F304AAE431F39FB265A188D08C6E3DF8E104603163F86490317",
    INIT_0d => x"A7A0A7A0A7FF8684A7A4A604263F8184A60A24C0DF8C21AEB9FE16480217068D",
    INIT_0e => x"E1FD0200CC1EE1FD0600CC393D3139F7265A0427A1ACA0A608C6E3DF8E1039A0",
    INIT_0f => x"178D0EE1FD20C60AE1FD08E1FD06E1FD5F04E1FD0100CC2E8D0CE1FDE000CC1E",
    INIT_10 => x"E1FCF92680C50EE1FC3B341F4AAF00C08EF42600C18C80E700E1FC218D00C08E",
    INIT_11 => x"54545454A6E6D0DF8E104444444462A6363439F92708C50EE1FC39F22740C50E",
    INIT_12 => x"FCBD8435FD265A20C60434B63562E762EA62A70F8462A65858585853A6E6E4E7",
    INIT_13 => x"0234A80117F12631813D273981230217F92653812A0217E2DF7F6802171186E3",
    INIT_14 => x"E0EB02340C2904358E01170434E46AE46AE4EBE0EBE0E6103421299101172629",
    INIT_15 => x"0117E26F1202161386E2DF731A02173F86BA27FFC102355FEB2080A70527E46A",
    INIT_16 => x"2320008310062762A3E4ECF901171286E3FCBDE4AF0130492562AC4D2930344A",
    INIT_17 => x"1780A684EB63EB62EB68011762AE750117981F03CB2F0017F3FE8E64E720C602",
    INIT_18 => x"10347120028D396532B701171486C326E4AC62AF5B0117981F53F526646A6501",
    INIT_19 => x"8D618D394AAF0229F68DF28D910017E50016F80016A101169035690017A4FE8E",
    INIT_1a => x"498D3944AF0229D58DD18D5E8D3946AF0229E08DDC8D728D3948AF0229EB8DE7",
    INIT_1b => x"8D3941A70229B18DB08D588D3942A70229BC8DBB8D6C8D3943A70229C78DC68D",
    INIT_1c => x"BF0016311FF48DB6FE8E39F726048180A63F011739C4A7808A0429A68DA58D5F",
    INIT_1d => x"8DC8FE8EE12044AED78DCEFE8EB4001643A6E18DD4FE8EF42048AEEA8DC2FE8E",
    INIT_1e => x"D02042A6B38DDFFE8ED92041A6BC8DDAFE8ECF204AAEC58DBCFE8ED82046AECE",
    INIT_1f => x"B2FE8EBF8DB88DB08DA98DA18D27FF17B2FE8E900016EBFE8EC4A6AA8DE4FE8E",
    INIT_20 => x"3C29088D011F42290E8DB800172D86121F4D29098DD520CE8DC78DC08D17FF17",
    INIT_21 => x"811D2530815B8D39E0AB04342829078D891F484848483229118D903561A71034",
    INIT_22 => x"3439021A39578003226681072561813937800322468112254181393080032239",
    INIT_23 => x"C602345120078B022F3981308B0F840235048D4444444402340235028D023510",
    INIT_24 => x"207F84048D0627E2DF7D00F09F6E8235F1265A3F8D438D2D860225E46880A608",
    INIT_25 => x"85E0DF9FA60234903501A6EE27018584A620E08E0926018584A6E0DFBE10342D",
    INIT_26 => x"3501A70235FA27028584A6E0DFBE1234458D2086008D8235018520E0B6052601",
    INIT_27 => x"A7FBDFFD0000CC30E08E39E2DFB7FF86016D84A7118684A70386E0DFBE138D90",
    INIT_28 => x"8D0427FEDF7D30E08E16345986028D1B86FEDF7F01E702C6FDDFFD04E703E702",
    INIT_29 => x"1A816C0027101B814100271008819635C5001784A70520098D042420810D2074",
    INIT_2a => x"51260A81110027100B812C0027100C81990027100D814500271016818E002710",
    INIT_2b => x"164A3327FBDFB67400165A3C0027105DFBDFFC9900168300261019C15CFBDFFC",
    INIT_2c => x"2710598116273DC1FEDFF65800160000CC5B00162500271050814CFBDFB66800",
    INIT_2d => x"2080FEDF7F39FDDFB70426FDDF7D39FEDF7F39FEDFB704263D81312754816E00",
    INIT_2e => x"A74C84E720C6FBDFB6168D0000CC1B20E12218C120C0FDDF7FFDDFF6ED224F81",
    INIT_2f => x"C15C4FF02650814CFBDFFC3903E702A7FBDFFDFCDFF64F39FEDF7FF726508102",
    INIT_30 => x"2650C15C84A702E7FBDFF72086FBDFF604E75F012519C15C04E6E78D5AEA2619",
    INIT_31 => x"FB0274FB0139FEDFF702E7FBDFF75FE4205F03E7FCDFF7082719C15CFCDFF6F4",
    INIT_32 => x"505EFA4CA5F847FDF8455CF94248FB1953FB183DFB1531FB105EFB047FFB0369",
    INIT_33 => x"94F9A7F8A7F8A7F8A7F894F992FC55D5F94488F958F1F853EDFB52A8F84DBCFA",
    INIT_34 => x"20205353455820524F4620342E312047554239305359530000000A0DFFFFFFFF",
    INIT_35 => x"43502020043D5053202004202D20043F54414857043E040000000A0D4B04202D",
    INIT_36 => x"20043D412020043D50442020043D58492020043D59492020043D53552020043D",
    INIT_37 => x"0000000000000000000004315343565A4E4948464504203A43432020043D4220",
    INIT_38 => x"300B2784AC1084AF1084EEAA558E10A0D08E84A7F086FB264A80A70F86F0FF8E",
    INIT_39 => x"2DA7D0DF8E10C0DFCE10FDFFB74444444443101F84EFD620ED26A0F08C00F089",
    INIT_3a => x"1084AF10AA558E1084EE2227A0F08C00F08930FB2A4AA66F0C862FA7F0862E6F",
    INIT_3b => x"2EA7D0DF8E10F186D520A5A70F88891F44444444101FD0DF8E1084EFE92684AC",
    INIT_3c => x"8EF32D0C814C80E7A66F0427A6E6211F4F2CE7A66F1420F92A4A0526A6E60C86",
    INIT_3d => x"9F6EC6DF9F6EC4DF9F6EC0DF9F6E62F816E2DFF753F9265A80A7A0A610C6F0FF",
    INIT_3e => x"0822CEDFBC8B300F27FFFF8CCCDFBE49584F4AAF80E64AAE431FCADF9F6EC8DF",
    INIT_3f => x"00FFB2FFC2FFBEFFBAFFB6FFC6FFB2FFC2DF9F6E42EE1F37F16E44AEC4EC1034"
    )

    port map (
	  do   => data_out1,
	  dop(0) => dp1,
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp1,
	  en   => cs1,
	  ssr  => rst,
	  we   => '0'
	);

my_mon : process ( rw, addr, cs, data_out0, data_out1 )
begin
    we    <= not rw;
	 cs0   <= '0';
    cs1   <= '0';
	 case addr(11) is
	 when '0' =>
	   cs0   <= cs;
		data_out <= data_out0;
    when '1' =>
		cs1   <= cs;
		data_out <= data_out1;
    when others =>
      null;
    end case;		
		
end process;

end architecture rtl;

