--===========================================================================--
--                                                                           --
--               Synthesizable PS/2 Keyboard Key map ROM for Spartan3        --
--                                                                           --
--===========================================================================--
--
--  File name      : keymap_rom2k_b16.vhd
--
--  Entity name    : keymap_rom 
--
--  Purpose        : Key code look up table for PS/2 Keyboard
--                   Converts 7 bit key code to ASCII
--                   Address bit 8      = Shift
--                   Address bit 7      = CAPS Lock
--                   Address bits 6 - 0 = Key code
--                   Data bits 6 - 0    = ASCII code
--                   Intended for Spartan 3/3E
--
--  Dependencies   : ieee.std_logic_1164
--                   ieee.std_logic_arith
--                   unisim.vcomponents
--
--  Uses           : RAMB16_S9
--
--  Author         : John E. Kent
--
--  Email          : dilbert57@opencores.org      
--
--  Web            : http://opencores.org/project,system09
--
--  Copyright (C) 2004 - 2010 John Kent
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--===========================================================================--
--                                                                           --
--                              Revision  History                            --
--                                                                           --
--===========================================================================--
--
-- Version Date        Author     Changes
--
-- 0.1     ????-??-??  John Kent  Initial version
-- 0.2     2010-06-17  John Kent  Revised Header, renamed data pins
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
library unisim;
	use unisim.vcomponents.all;

entity keymap_rom is
    Port (
       clk      : in  std_logic;
       rst      : in  std_logic;
       cs       : in  std_logic;
       rw       : in  std_logic;
       addr     : in  std_logic_vector (8 downto 0);
       data_in  : in  std_logic_vector (7 downto 0);
       data_out : out std_logic_vector (7 downto 0)
    );
end keymap_rom;

architecture rtl of keymap_rom is


signal we : std_logic;
signal dp : std_logic;
signal ad : std_logic_vector(10 downto 0);

begin

  ROM : RAMB16_S9
    generic map (
    INIT_00 => x"00327761737a0000003171000000000000600900000000000000000000000000",
    INIT_01 => x"003837756a6d00000036796768626e0000357274667620000033346564786300",
    INIT_02 => x"00005c005d0d000000003d5b00270000002d703b6c2f2e000039306f696b2c00",
    INIT_03 => x"0000000000000000001b000000007f0000000000000000000008000000000000",
    INIT_04 => x"00121701131a0000001111000000000000000900000000000000000000000000",
    INIT_05 => x"001817150a0d00000016190708020e0000151214061600000013140504180300",
    INIT_06 => x"00001c001d0d000000001d1b00070000000d101b0c0f0e000019100f090b0c00",
    INIT_07 => x"0000000000000000001b000000001f0000000000000000000008000000000000",
    INIT_08 => x"00405741535a00000021510000000000007e0900000000000000000000000000",
    INIT_09 => x"002a26554a4d0000005e594748424e0000255254465620000023244544584300",
    INIT_0A => x"00007c007d0d000000002b7b00220000005f503a4c3f3e000028294f494b3c00",
    INIT_0B => x"0000000000000000001b000000007f0000000000000000000008000000000000",
    INIT_0C => x"00001701131a00000001110000000000001e0900000000000000000000000000",
    INIT_0D => x"000a06150a0d0000001e190708020e0000051214061600000003040504180300",
    INIT_0E => x"00001c001d0d000000001d1b00020000001f101a0c1f1e000008090f090b1c00",
    INIT_0F => x"0000000000000000001b000000001f0000000000000000000008000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do     => data_out,
	  dop(0) => dp,
	  addr   => ad,
	  clk    => clk,
	  di     => data_in,
	  dip(0) => dp,
	  en     => cs,
	  ssr    => rst,
	  we     => we
	);

my_keymap_rom_b16 : process ( rw, addr )
begin
	 we    <= not rw;
    ad(8 downto 0) = addr;
    ad(10 downto 9) = "00";
end process;

end architecture rtl;

