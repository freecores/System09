sys09bug_rom_inst : sys09bug_rom PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
