-- $Id: Maisforth_rom16k_b16.vhd,v 1.2 2008-03-14 15:52:43 dilbert57 Exp $
--===================================================================
--
-- Mais Forth 16K ROM for the 6809 
-- Made from Block RAM
--	Resides from C000 to 3FFF
-- with I/O at $B000 to $B0FF
-- (6850 ACIA at $B000)
-- (PS/2 Keyboard at $B010)
-- (VDU8 at $B020)
--
--===================================================================
--
-- Date: 24th April 2006
-- Author: John Kent
--
-- Revision History:
-- 24 April 2006 John Kent
-- Initial release
--
-- 29th June 2005 John Kent
-- Added CS term to CE decodes.
--
-- 10th August 2007 John Kent
-- Turned into 16K Byte Mais Forth ROM.
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
library unisim;
	use unisim.vcomponents.all;

entity maisforth_rom_16k is
    Port (
       clk   : in  std_logic;
		 rst   : in  std_logic;
		 cs    : in  std_logic;
		 rw    : in  std_logic;
       addr  : in  std_logic_vector (13 downto 0);
       rdata : out std_logic_vector (7 downto 0);
       wdata : in  std_logic_vector (7 downto 0)
    );
end maisforth_rom_16k;

architecture rtl of maisforth_rom_16k is


signal we    : std_logic;
signal dp    : std_logic_vector(7 downto 0);
signal ce    : std_logic_vector(7 downto 0);
signal rdata_0 : std_logic_vector(7 downto 0);
signal rdata_1 : std_logic_vector(7 downto 0);
signal rdata_2 : std_logic_vector(7 downto 0);
signal rdata_3 : std_logic_vector(7 downto 0);
signal rdata_4 : std_logic_vector(7 downto 0);
signal rdata_5 : std_logic_vector(7 downto 0);
signal rdata_6 : std_logic_vector(7 downto 0);
signal rdata_7 : std_logic_vector(7 downto 0);

begin

  RAM0 : RAMB16_S9
    generic map ( 
    INIT_00 => x"F9E8FAB4FBDDFB0CFABAFA15FBCEFAA5FAE9F7A5F7FEFA7BFADFF8F0F85EF17E",
    INIT_01 => x"00000200000000000000003000F3FB1F000000000003037AEA0FFDC1ED63FA61",
    INIT_02 => x"003B00003B00003B00003B00000A000000000000000003000003000000000000",
    INIT_03 => x"20375449584504020000846E0635011F45545543455845070200003B00003B00",
    INIT_04 => x"0000B16E20370227063500008310455552542D4E4F2D544958450C040000B16E",
    INIT_05 => x"4404040000B16E2037022606350000831045534C41462D4E4F2D544958450D04",
    INIT_06 => x"6E101F063410352035203653454F444F4406040000B16E10362037211F455649",
    INIT_07 => x"36EEC0BD3A4F44030400007EC03DCDD5C0BDEEC0BD52454F444F4406040000B1",
    INIT_08 => x"05040000B16E101F06341035EEC0BD4554414552434F440804BEC0B16E203520",
    INIT_09 => x"341035EEC0BD4E4F43434F4406040000B16E101F06341035EEC0BD5241564F44",
    INIT_0a => x"4F440504E4C0B16E84EC06341035EEC0BD4E4F434F440504F8C0B16E1D84E606",
    INIT_0b => x"EC06341035EEC0BD524156494F4406045DC1B16E84EC06341035EEC0BD4C4156",
    INIT_0c => x"41564F440604CEC0B16E94EC06341035EEC0BD4C4156494F4406041FC1B16E84",
    INIT_0d => x"1D5A012702845F00B0B606343F54494D45050285C0B16EE1E34958EEC0BD5352",
    INIT_0e => x"552106060000B16E063501E7FA27028484A600B08E54494D4528050486C1B16E",
    INIT_0f => x"2701845F00B0B606343F59454B04020000B16E063584A7558600B08E54524153",
    INIT_10 => x"070468C0B16E4F01E6FA2701C484E600B08E063459454B0302F2C1B16E1D5A01",
    INIT_11 => x"C4AE063424454E494C4E49070479C0B16EC4AF81ECC4AE063423454E494C4E49",
    INIT_12 => x"C4AF853080E6C4AE063424454E494C4E492F08040000B16EC4AF3A10344F80E6",
    INIT_13 => x"3500008310292846490404A1C0B16EA4AE1029284F544F47060434C2B16E0635",
    INIT_14 => x"052706350000831029284F52455A4649080476C2B16E2231B16EA4AE10052606",
    INIT_15 => x"A0E6063429432803040000B16EA1EC0634292802040000B16E2231B16EA4AE10",
    INIT_16 => x"84E3A1AE29284F542B050467C2B16E063584EDA1AE29284F540404B8C2B16E1D",
    INIT_17 => x"C2B16E063584ED0100C384EC0634A1AE292852434E4906041FC2B16E063584ED",
    INIT_18 => x"05040000B16E063510368B300636E1A30080CC011F1036A1AE29284F440404C6",
    INIT_19 => x"EC06342928504F4F4C060402C3B16EA4AE1006356232DD26E4A31029284F443F",
    INIT_1a => x"504F4F4C2B070408C2B16E063546332231B16EA4AE100635C4ED09290100C3C4",
    INIT_1b => x"33504F4F4C4E550602D6C2B16E20374433455641454C0502ACC2DE20C4E32928",
    INIT_1c => x"0493C3B16E48A346EC06344A01029BC1B16E42A3C4EC0634490102AEC1B16E46",
    INIT_1d => x"54060449C1250090C1BD47534D504F54060469C3230090C1BD434F56504F5406",
    INIT_1e => x"444C480304BEC3290090C1BD41464E504F54060408C1270090C1BD584650504F",
    INIT_1f => x"0090C1BD23534303041FC32D0090C1BD545845544E4F4307044DC22B0090C1BD",
    INIT_20 => x"04E9C2330090C1BD45444F4D0404E8C3310090C1BD322D2347534D0604DDC12F",
    INIT_21 => x"03048FC2370090C1BD53454D495423060478C3350090C1BD4E4F495443455307",
    INIT_22 => x"0090C1BD45524548540504A0C33B0090C1BD424902045AC3390090C1BD424923",
    INIT_23 => x"4D4948050636C3410090C1BD5245560306CDC33F0090C1BD524F48030633C13D",
    INIT_24 => x"C3470090C1BD3F544F44040656C4450090C1BD4B4F020604C4430090C1BD4D45",
    INIT_25 => x"BD4E493E030270C44B007BC1BD445257030420C4490090C1BD455245480402AF",
    INIT_26 => x"C453007BC1BD4554415453050230C451007BC1BD45534142040271C14F007BC1",
    INIT_27 => x"2705068AC458007BC1BD3249575327050613C455007BC1BD334957532705064B",
    INIT_28 => x"C1BD4957532704060CC55E007BC1BD515249270406E2C45B007BC1BD51524946",
    INIT_29 => x"C100C052C1BD4E494749524F06023FC464007BC1BD494D4E27040619C561007B",
    INIT_2a => x"C37F3DC1BD544E45525255430704F0C4753DC1BD4B43415453444E49460904C5",
    INIT_2b => x"0152C1BD3052020495C47E0152C1BD3053020433C5800052C1BD4249540304DC",
    INIT_2c => x"070484C5FC0252C1BD305343030486C3000252C1BD465542594C460604A2C4FE",
    INIT_2d => x"BD455552540402BBC4023DC1BD4C4C454304066EC57E3DC1BD455A4953424954",
    INIT_2e => x"4C430704F8C3203DC1BD4C4202029FC5003DC1BD45534C41460502C7C4FF3DC1",
    INIT_2f => x"0493C5B16EFE01CE522D5241454C430704AEC5B16E06357E01CE10532D524145",
    INIT_30 => x"35011F21430202DDC5B16E301F06344050520304BAC5B16E401F063440505303",
    INIT_31 => x"0635011F21320202C6C5B16E063584ED0635011F21010253C5B16E063584E706",
    INIT_32 => x"0306D4C4B16E063584ED84E30635011F212B0202FEC4B16E063584ED063581ED",
    INIT_33 => x"3584ED0100C384EC011F212B31030600C6B16E063584E784EB0635011F212B43",
    INIT_34 => x"32020279C5B16E84EC011F40010242C5B16E4F84E6011F40430202F0C5B16E06",
    INIT_35 => x"060DC6B16E10344F80E6011F544E554F43050272C6B16E103484AE81EC011F40",
    INIT_36 => x"3706343E5202027CC4B16E06350636523E0202D3C5B16E103481EC011F2B4002",
    INIT_37 => x"37063706343E52320302CEC6B16E0635063610361035523E3203029EC6B16E06",
    INIT_38 => x"C4EC103442AE06344052320302C0C6B16EC4EC063440520202E6C6B16E103410",
    INIT_39 => x"0225C7B16E4433504F52445232060608C7B16E4233504F5244520506DAC6B16E",
    INIT_3a => x"04024FC7B16E10340634E4AE505544320402F7C6B16E06356232504F52443205",
    INIT_3b => x"C7B16E66EC063466EC06345245564F3205025FC7B16E10346432103550494E32",
    INIT_3c => x"5432050264C4B16E62AF62EC1037E4ED64AF64ECE4AE06365041575332050240",
    INIT_3d => x"C088C7FBC688C7EAC6FFC0BD544F5232040232C77EC075C788C7FFC0BD4B4355",
    INIT_3e => x"C6B16E0635504F5244040293C6B16E06340227000083105055443F0402AEC67E",
    INIT_3f => x"504157530402AFC4B16E62EC06345245564F040286C6B16E0634505544030239"
    )

    port map (
	  do   => rdata_0,
	  dop(0) => dp(0),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => wdata,
	  dip(0) => dp(0),
	  en   => ce(0),
	  ssr  => rst,
	  we   => we
	);

  RAM1 : RAMB16_S9
    generic map (
	 INIT_00 => x"AE544F52030282C7B16E1034E4EDE4AE4B43555404026FC7B16E101FE4EDE4AE",
    INIT_01 => x"4E03020BC8B16EE4AFE4EC62ED62AE544F522D040226C5B16E62AF62ECE4EDE4",
    INIT_02 => x"E4A3104E494D03025FC6B16E84EC3A411F584B43495004021BC8B16E62325049",
    INIT_03 => x"A3104E494D5504061AC6B16E0635D02EE4A31058414D03024DC6B16E0635E02D",
    INIT_04 => x"891F3C3002029DC7B16E0635AE22E4A31058414D5504062CC8B16E0635BF25E4",
    INIT_05 => x"103E300202D6C7B16E5F4FB16E1D530426000083103D3002023EC8B16E891F1D",
    INIT_06 => x"0202E2C7B16E5F4FD927E1A33D0102FBC7B16E891F431D891FB16E0226000083",
    INIT_07 => x"3E55020269C8B16EEE26000083103E3C3003029BC8B16EFFFFCC0327E1A33E3C",
    INIT_08 => x"4FC72DE1A33E010249C8B16E5F4FD422E1A33C5502028AC8B16E5F4FE225E1A3",
    INIT_09 => x"02D2C8B16EE0E4E0A4444E4103020BC9B16E5F4FBA2EE1A33C0102EEC8B16E5F",
    INIT_0a => x"545245564E49060279C8B16EE0E8E0A8524F58030226C9B16EE0EAE0AA524F02",
    INIT_0b => x"A8C8B16EFA261F304958062784300635011F54464948534C060262C5B16E5343",
    INIT_0c => x"45545942080681C9B16EFA261F305644062784300635011F5446494853520602",
    INIT_0d => x"14C7B16E0100832D31020240C9B16E0100C32B310202C4C7B16E891E50415753",
    INIT_0e => x"2D0102B6C9B16EE1E32B010259C9B16E56472F320202BCC8B16E49582A320202",
    INIT_0f => x"19C9B16E4959101F063449580635011F2A3244030267C9B16E0100C35343E1A3",
    INIT_10 => x"B16EE820442F3255440406AFC7B16E101F063456460635011F56472F32440302",
    INIT_11 => x"06D5C9B16EEF2D4D5342410302EDC7B16E0100C3534345544147454E0602ECC9",
    INIT_12 => x"011F1D5F063445544147454E4407029BC9B16EDD2D06354D45544147454E3F07",
    INIT_13 => x"443F080633C9B16EE22D4D53424144040252CAB16EE1A31D00C2101F62ED62A3",
    INIT_14 => x"8900C9101F62ED62E30635011F2B44020216CAB16ECF2D06354D45544147454E",
    INIT_15 => x"C9B16E6632E4A3008200C264EC66ED62A366EC06342D44020201CAB16EE1E300",
    INIT_16 => x"ED3D61E665A616342A4D55030259C8B16E008900C9063562ED62E32B4D0202DE",
    INIT_17 => x"E33D64A6E4A7E4E649008661ED61E33DE4E665A661ED008962EB3D61E664A662",
    INIT_18 => x"626963696469656810008E0634444F4D2F4D5506027DCAB16EE4AF643262AEE4",
    INIT_19 => x"62AE534364ECE2261F306469656962ED0225E4A30620FE1C62EDE4A3082462EC",
    INIT_1a => x"370635FA261F30A0E7062700008C303520364C4C49460402C1C9B16E643264AF",
    INIT_1b => x"C20927A0A080A60F205FE4EDE4AE1062AF1062AE62E33E3C530306C2CAB16E20",
    INIT_1c => x"AF1062AE62E345564F4D430502D4CAB16E30351DED26E4ACB16E303501CA1D00",
    INIT_1d => x"3E45564F4D4306022AC6B16E06353035F826E4ACA0E780E60420E4EDE4AE1062",
    INIT_1e => x"343F31B16E06353035F726E4AC10A2E782E60420AB31E4AE1062AF108B3062AE",
    INIT_1f => x"F8261F30E126A0E1082700008C3035203650494B53040666CBB16E101F203720",
    INIT_20 => x"02FDC8C220F8261F30C627A0E1082700008C303520364E4143530406ABC9DD20",
    INIT_21 => x"4F423E0502DFC8B16E0100C32B52414843050220CCB16E0200C32B4C4C454305",
    INIT_22 => x"00832D5241484305064ACCB16E0200832D4C4C4543050694CBB16E0300C35944",
    INIT_23 => x"74CCB16E4958534C4C454305022ECCB16E0300833E59444F42050690CAB16E01",
    INIT_24 => x"52040266CCB16E0300834B4E494C3E454D414E090423CAB16E53524148430503",
    INIT_25 => x"CBC97EC0DBC7C0CB7ACCAEC9DDC626CCE6C704C64EC80BC7D1C6FFC0BD4C4C4F",
    INIT_26 => x"00DCC2FFC0BD544F4C4C41050258CC7EC0D7C940BCC2A7C4FFC0BD4441500302",
    INIT_27 => x"FFC0BD2C430202EACB7EC04900DCC2B3C52CC6A7C4FFC0BD2C01024CC97EC049",
    INIT_28 => x"CCB16E101F85301FC480E6011F3E454D414E0506A8CA7EC04900F0C21DC6A7C4",
    INIT_29 => x"FFC0BD52454F4421050481CCB16E101FFA2682E460C6011F454D414E3E0506E6",
    INIT_2a => x"040DCDB16E1D5A5801C482E6011F4D4D494004049ECC7EC02CC6AEC913CDD4C3",
    INIT_2b => x"CCB16E1D7EC482E6011F434F5640040460CDB16E891F1D82E6011F3F4D4F4804",
    INIT_2c => x"0405CCB16E1D5A012400C6E1A3E4AFE1A362EC011FE4A34E49485449570602FA",
    INIT_2d => x"BD53433E0304C1CC7EC0E0C937C97CBCC2C4C97ACCFCC397C5FFC0BD50534303",
    INIT_2e => x"00DCC2FFBCC2A1C6A4CDFFC0BD3E5343030482CD7EC03CC6A4CD2F00F0C2FFC0",
    INIT_2f => x"C2DDC6D3CD2F00DCC22ACAD1C6FCC3FFC0BD4B4349502D5343070240CA7EC02F",
    INIT_30 => x"26CE25C300BCC20BC7D1C6FFC0BD4C4C4F522D53430702B9CB7EC0BFCD2F00CB",
    INIT_31 => x"CE7EC0BFCDFBC633CE3DC3BFCD39CE25C300BCC2EAC6D3CDDDC620CE3DC3D3CD",
    INIT_32 => x"38CAF2C738CAF2C7FFC0BD2A4D020237CDB16E891F1D891F0634443E5303020A",
    INIT_33 => x"C775CAD1C6D1C6F2C7FFC0BD4D45522F4D53060252CE7EC086CA50C988C7D8CA",
    INIT_34 => x"4F4D2F4D46060271CD7EC000C848CADDC600C848CA50C90BC7DDC613CB38CA0B",
    INIT_35 => x"9EC850C90BC71FC800C848CA0BC700C813CB38CA0BC775CA10C8D1C6FFC0BD44",
    INIT_36 => x"BD2A01024DCD7EC02BC700C8E0C91FC80BC7B9C9D6CE7BC2F2C72ACAD6CE7BC2",
    INIT_37 => x"020CCB7EC0A1CEDDC646CED1C6FFC0BD444F4D2F040242CE7EC0DBC755CEFFC0",
    INIT_38 => x"2A05029ACE7EC0DBC7F0CEFFC0BD444F4D0302E6CD7EC042C8F0CEFFC0BD2F01",
    INIT_39 => x"7EC042C824CFFFC0BD2F2A02028CCC7EC0A1CEDDC655CED1C6FFC0BD444F4D2F",
    INIT_3a => x"C10DBCC2FFC0BD52430202A0CD7EC03F00F0C2CBC1FFC0BD54494D450402D4CC",
    INIT_3b => x"D6C5FFC0BD4543415053050243CF7EC04100F0C23F00CBC2CCC5CBC10ABCC2CB",
    INIT_3c => x"48CFE6C7A4CF25C300BCC200C8D6C5FFC0BD534543415053060275CF7EC048CF",
    INIT_3d => x"3DC348CFB4C6C2CF25C300BCC2FFC0BD45505954040249CB7EC0DBC79CCF3DC3",
    INIT_3e => x"CBC2CCC53F00CBC2CCC548CF0CBCC2FFC0BD454741500402DDCE7EC0DBC7BACF",
    INIT_3f => x"C1F2C7D6C508BCC2AFC068C4FFC0BD45434150534B434142090634CF7EC04100" 
    )

    port map (
	  do   => rdata_1,
	  dop(0) => dp(1),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => wdata,
	  dip(0) => dp(1),
	  en   => ce(1),
	  ssr  => rst,
	  we   => we
	);

  RAM2 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0CC2FFC0BD474E49545045434341090434CA7EC03F00DCC2FFBCC2CBC1CBC1CB",
    INIT_01 => x"D4C808BCC27EC0DBC764C73BD07BC2D4C8F2C70DBCC254D07BC228C9D6C5E6C7",
    INIT_02 => x"D07BC2D4C84EC804BCC2F2C7D6C51ED06EC2B9C9F1CF4ED07BC2E6C752D07BC2",
    INIT_03 => x"504543434106026DCE1ED06EC2AEC948CF1DC6D7C975C7E6C71ED06EC2DBC767",
    INIT_04 => x"CB00C8CCC510C8FFC0BD444F4D2F55440606BBCD7EC01BD0CCC500C8FFC0BD54",
    INIT_05 => x"C6D8CAD1C6DBC7D8CA10C8FFC0BD2A55440306E7CF7EC0DDC613CB00C8D1C613",
    INIT_06 => x"0270CA7EC01DC6E0C32B00DCC2FFBCC2FFC0BD444C4F48040222CD7EC0D7C9DD",
    INIT_07 => x"09BCC2E6C7FFC0BD54494749443E0604ABCF7EC02B00CBC2C5CCFFC0BD233C02",
    INIT_08 => x"1FC896D095C6CCC4FFC0BD2301027AD07EC0D7C930BCC2D7C937C907BCC21BC9",
    INIT_09 => x"230202EBCE7EC02FD198C243C954C715D1FFC0BD5323020287CF7EC0CDD0F8D0",
    INIT_0a => x"C2AFC09EC8FFC0BD4E474953040256CF7EC0E0C9F2C7C5CCE0C346C7FFC0BD3E",
    INIT_0b => x"C9CF7EC041D12CD1E3D0FFC0BD474E495254532E55440906F1D07EC0CDD02DBC",
    INIT_0c => x"06AED07EC041D158D11FC82CD1E3D075CA10C8FFC0BD474E495254532E440806",
    INIT_0d => x"D1FFC0BD2E554403068FD07EC0B0CF8ECFE0C95DC854C7FFC0BD455059545205",
    INIT_0e => x"0202CAD17EC0A6D1DDC673D1D1C6FFC0BD522E55440406C8D07EC07BCFB0CF73",
    INIT_0f => x"021ECF7EC0BCD100BCC2FFC0BD2E55020213D17EC07BCFB0CF8AD1FFC0BD2E44",
    INIT_10 => x"D17EC0A6D1DDC68AD1D1C6FFC0BD522E440302A0D17EC0E2D146CEFFC0BD2E01",
    INIT_11 => x"C6FFC0BD522E0202E0D07EC0A6D1DDC673D100BCC2D1C6FFC0BD522E55030229",
    INIT_12 => x"4345440702DFD17EC002D295C6FFC0BD3F010200CF7EC0A6D1DDC68AD146CED1",
    INIT_13 => x"C6CCC410BCC2FFC0BD5845480302B8D17EC02CC6CCC40ABCC2FFC0BD4C414D49",
    INIT_14 => x"554F530602F0D17EC02CC6CCC402BCC2FFC0BD5952414E494206063CCC7EC02C",
    INIT_15 => x"AFE4EC62ED62E3011F474E495254532F070222D27EC043C44EC4FFC0BD454352",
    INIT_16 => x"435441432906049CD2B16E10365E304036284843544143060411D0B16EE1A3E4",
    INIT_17 => x"0469D17EC0E1D270C0CFD2FFC0BD484354414305023ED1B16E5F4F0634443348",
    INIT_18 => x"524F42410502AFD2B16E2037101F4037F926C1A310301F011F574F5248542806",
    INIT_19 => x"6E20C002227AC1062561C1524550505528060473D27EC007D3FFBCC2FFC0BD54",
    INIT_1a => x"AEC91DC6F2C735D389C6E6C764D325C300BCC2FFC0BD524550505505064ED2B1",
    INIT_1b => x"7EC8D1C6E0C954C71FC8FFC0BD455241504D4F43070244D37EC0DBC754D33DC3",
    INIT_1c => x"4F4D0402ECD27EC0AEC9C4C9BFC8AFC0E6C7DDC67EC02BC78CD37BC2C9C76ACB",
    INIT_1d => x"414C50050600D37EC0C0CB7EC09ACBB5D37BC289CD75C7D7C954C7FFC0BD4556",
    INIT_1e => x"A3D2D1C6FFC0BD44524F57040253D17EC0A2D300C834CC1DC654C7FFC0BD4543",
    INIT_1f => x"3CC6B3C454C7E0C9F2C7D1C60ACCDDC600C8F2C7EFCB0BC710C8B7D295C6BFC4",
    INIT_20 => x"BD45535241500502BCD37EC0A7C450C6BFC4E0C9D7C9F2C8E6C7DDC6C2D3A7C4",
    INIT_21 => x"BFC4E0C9D7C9F2C8E6C7DDC6EAC60ACCDDC654C7B7D295C6BFC4A3D2D1C6FFC0",
    INIT_22 => x"C6B16E0635042B5D401F06344B434154533F0606DAD27EC0E0C9F2C7DDC650C6",
    INIT_23 => x"CD49BCC202BCC295C6CCC4FFC0BD455341423F05064DD407D37E1D5C01264DFC",
    INIT_24 => x"D3EABCC292C0D4C8FFC0BD524941503F0506D4D37EC007D3C2BCC264D292C089",
    INIT_25 => x"0802A6D47EC007D3F2BCC292C095C6DAC4FFC0BD504D4F433F0506C8D27EC007",
    INIT_26 => x"4D4F4309046BD37EC04900DCC2B3C52CC6A7C4ACD4FFC0BD2C454C49504D4F43",
    INIT_27 => x"CD7EC02CC6DAC4CCC5FFC0BD5B01030ECF7EC0C8D427C2FFC0BD2928454C4950",
    INIT_28 => x"FFC0BD45524548542D454641530A046CD47EC02CC6DAC4BFC5FFC0BD5D0102CF",
    INIT_29 => x"594C46050400D27EC05CC43D00CBC28BC535D57BC20EC9E0C98BC55CC440BCC2",
    INIT_2a => x"C004D5EAC6DDC64900CBC2E6C73D00CBC2A7C41DD592C095C6DAC4FFC0BD5245",
    INIT_2b => x"FFC0BD2953282204045CD27EC03D00CBC24900CBC25CC4A7C4F4D47EC0E6D4C3",
    INIT_2c => x"C2FFC0BD282E02033CD57EC0B0CF3CC2FFC0BD295328222E050486D27EC03CC2",
    INIT_2d => x"78D57EC0DACCAEC989C6D9D3FFC0BD2C44524F570506BFD47EC0B0CF1FD429BC",
    INIT_2e => x"4F424109049DD37EC0C2D3DACCAEC9F2C7A7C41FD4FFC0BD2C45535241500606",
    INIT_2f => x"06031BD37EC056C207D3FEBCC23100CBC20BC7F8D57BC2FFC0BD295328225452",
    INIT_30 => x"42D5FFC0BD22010739D27EC0C8D522BCC2E6D5E6D442D5FFC0BD2254524F4241",
    INIT_31 => x"42D5FFC0BD222E020319D61ED66EC2FFC0BD225302038FD40FD66EC27DD5E6D4",
    INIT_32 => x"00CBC2E8CCB6C3E8CC00C8A7C4FFC0BD2247534D0406F2D40FD66EC28DD5E6D4",
    INIT_33 => x"0438D67EC0CEC9E0C900C871C504C6FFC0BD48545045440502C1D50FD66EC225",
    INIT_34 => x"45444F4D54494E49080402D57EC089CD8000AFC280BCC2FFC0BD3F5449423805",
    INIT_35 => x"C1BCC2AFC0FFC0BD4C4147454C4C493F0804DCD57EC03300CBC230BCC2FFC0BD",
    INIT_36 => x"BCC2B9C900C83300CBC220BCC2FFC0BD4745525845444E490804AFD67EC007D3",
    INIT_37 => x"BCC2FFC0BD45444F4347455207042ED37EC043C96EC905BCC2B8D60EC9F2C703",
    INIT_38 => x"4040201006040200535559584442412C107DD5D1C6E0C937C9D6C528C9F2C75A",
    INIT_39 => x"45444F4D2B0504DCD407D3C1BCC27EC089C6D7C932D77BC20ACCDDC610C8CEC9",
    INIT_3a => x"040ED27EC037C90FBCC292C0E2C850BCC237C9F000AFC2E6C7D7C918C4FFC0BD",
    INIT_3b => x"AFC200C88AD77BC286D6E6C7E0C9D7C902BCC2A7C400C8FFC0BD4C4552435005",
    INIT_3c => x"C0BD544553464F43060497D67EC0E8CCFDCC00C8B9C97EC0FDCCFDCC37C9FE00",
    INIT_3d => x"10BCC2F0BCC2F2C77EC0DBC7FDCC43C904BCC237C9F000AFC2B8D798C2F2C7FF",
    INIT_3e => x"CC43C937C91FBCC200C837C960BCC2E3D77BC237C9ABC837C910BCC2F2C789CD",
    INIT_3f => x"04FFD57EC0E8CCFDCC7EC0FDCCFDCC37C9FE00AFC2F7D77BC286D6F2C77EC0FD"
    )

    port map (
	  do   => rdata_2,
	  dop(0) => dp(2),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => wdata,
	  dip(0) => dp(2),
	  en   => ce(2),
	  ssr  => rst,
	  we   => we
	);

  RAM3 : RAMB16_S9
    generic map ( 
    INIT_00 => x"C725D87BC2D4C88900AFC2E6C737C98F00AFC2E6C7FFC0BD44455845444E4907",
    INIT_01 => x"C2D4C88F00AFC2E6C77EC066D7DBC737D87BC2D4C88D00AFC2E6C77EC09ED7DB",
    INIT_02 => x"C989C6FFC0BD44454D4D4905043AD77EC0FDCCDBC77EC0E8CCFDCCDBC74BD87B",
    INIT_03 => x"D5C0BDEEC0BD5845534F44050468D67EC0FDCC7EC0E8CC6DD87BC2B8D646CEB9",
    INIT_04 => x"7EC0A0D6E8CC95C6D5C0BDEEC0BD324957534F44060487D57EC0A0D6FDCC89C6",
    INIT_05 => x"ABD57EC0A0D6FDCCFDCC89C6B8D618C4D5C0BDEEC0BD494157434F44060419D4",
    INIT_06 => x"7EC05AD8DBC7E0D87BC2D4C800BCC2E6C7A0D618C4FFC0BD5244414E45470604",
    INIT_07 => x"DBC706D97BC2D4C820BCC2E6C77EC0FDCCDBC7DBC7F3D87BC2D4C810BCC2E6C7",
    INIT_08 => x"04A3D87EC0B8D67EC0E8CCDBC7DBC719D97BC2D4C830BCC2E6C77EC008D8DBC7",
    INIT_09 => x"BD59444C4F44050480D67EC0C8D8FDCC40D7B4C6D5C0BDEEC0BD47454E4F4405",
    INIT_0a => x"89C6D5C0BDEEC0BD4758454F44050420D97EC0C8D8E8CC40D7C3C6D5C0BDEEC0",
    INIT_0b => x"D5C0BDEEC0BD41454C4F44050439D97EC0A0D6FDCCD7C96EC904BCC200C8FDCC",
    INIT_0c => x"BDEEC0BD5145424F44050474D97EC0A0D608D8FDCC89C6B8D6E0C920BCC218C4",
    INIT_0d => x"C0FDCCFDCC00C8C1D97BC286D6E6C7A0D6E0C9D7C902BCC2A7C400C889C6D5C0",
    INIT_0e => x"BDEEC0BD4152424F44050496D97EC0E8CCE0C902BCC2FDCC00C8FDCC10BCC27E",
    INIT_0f => x"CCFDCCA4C900C803DA7BC286D6E6C7A0D6E0C9D7C902BCC2A7C400C895C6D5C0",
    INIT_10 => x"C0D0D689C6D5C0BDEEC0BD292D4F44040499D57EC0E8CCB9C9FDCC00C87EC0FD",
    INIT_11 => x"52534C0308F3D6004329D9BD4D4F43030854D8004029D9BD47454E030860D77E",
    INIT_12 => x"0830DA004729D9BD52534103084BD6004629D9BD524F52030881D1004429D9BD",
    INIT_13 => x"4929D9BD4C4F52030810DA004829D9BD4C534C03088BD8004829D9BD4C534103",
    INIT_14 => x"545354030874D8004C29D9BD434E49030897D7004A29D9BD434544030852D900",
    INIT_15 => x"0812D5004F29D9BD524C430308C1D8004E29D9BD504D4A030878DA004D29D9BD",
    INIT_16 => x"BD414342530408CDDA018129D9BD41504D430408C0DA018029D9BD4142555304",
    INIT_17 => x"9CDA018429D9BD41444E41040890DA028329D9BD444255530408B4DA018229D9",
    INIT_18 => x"D9BD415453030800D8018629D9BD41444C0308D6D9018529D9BD415449420408",
    INIT_19 => x"08DADA018929D9BD414344410408F4DA018829D9BD41524F450408C7D6008729",
    INIT_1a => x"D9BD58504D4304084CDB018B29D9BD41444441040833DB018A29D9BD41524F03",
    INIT_1b => x"5303082BD6028E29D9BD58444C030801DB008D29D9BD52534A03080EDB028C29",
    INIT_1c => x"C129D9BD42504D4304088ADB01C029D9BD42425553040826DB008F29D9BD5854",
    INIT_1d => x"41040860DA02C329D9BD44444441040854DA01C229D9BD42434253040897DB01",
    INIT_1e => x"C629D9BD42444C03083CDA01C529D9BD425449420408A8DA01C429D9BD42444E",
    INIT_1f => x"44410408BEDB01C829D9BD42524F45040840DB00C729D9BD4254530308E7DA01",
    INIT_20 => x"01CB29D9BD424444410408FDDB01CA29D9BD42524F0308A4DB01C929D9BD4243",
    INIT_21 => x"BD55444C030848DA00CD29D9BD44545303080ADC02CC29D9BD44444C03086CDA",
    INIT_22 => x"F0DB02831042D9BD44504D430408E4DB00CF29D9BD555453030816DC02CE29D9",
    INIT_23 => x"59545303081ADB028E1042D9BD59444C030866DB028C1042D9BD59504D430408",
    INIT_24 => x"00CF1042D9BD5354530308B1DB02CE1042D9BD53444C0308CBDB008F1042D9BD",
    INIT_25 => x"040824DA028C1142D9BD53504D43040847DC02831142D9BD55504D43040896DC",
    INIT_26 => x"327DD9BD5341454C04083BDC317DD9BD5941454C040884DA307DD9BD5841454C",
    INIT_27 => x"D9BD5246540308BFDC1E5BD9BD47584503082FDC337DD9BD5541454C040889DC",
    INIT_28 => x"4141440308D7DC137DD8BD434E59530408B1DC127DD8BD504F4E03086FDC1F5B",
    INIT_29 => x"424103087CDC397DD8BD535452030823DC1D7DD8BD58455303087EDB197DD8BD",
    INIT_2a => x"5303083DDD3D7DD8BD4C554D0308A3DC3B7DD8BD4954520308FADC3A7DD8BD58",
    INIT_2b => x"CBDC437DD8BD414D4F43040861DC407DD8BD4147454E040848DD3F7DD8BD4957",
    INIT_2c => x"D8BD41525341040859DB467DD8BD41524F52040872DB447DD8BD4152534C0408",
    INIT_2d => x"4F5204088DDD487DD8BD414C534C040881DD487DD8BD414C5341040899DD477D",
    INIT_2e => x"C9DD4C7DD8BD41434E49040853DC4A7DD8BD414345440408E3DC497DD8BD414C",
    INIT_2f => x"D8BD4247454E04081CDD4F7DD8BD41524C43040875DD4D7DD8BD415453540408",
    INIT_30 => x"4F520408E1DD547DD8BD4252534C040832DD537DD8BD424D4F430408EFDC507D",
    INIT_31 => x"11DE587DD8BD424C5341040829DE577DD8BD42525341040810DD567DD8BD4252",
    INIT_32 => x"D8BD424345440408BDDD597DD8BD424C4F5204081DDE587DD8BD424C534C0408",
    INIT_33 => x"4C43040805DE5D7DD8BD42545354040859DE5C7DD8BD42434E4904085EDD5A7D",
    INIT_34 => x"3F1195D8BD33495753040835DE3F1095D8BD3249575304087DDE5F7DD8BD4252",
    INIT_35 => x"48535004084DDE1CADD8BD4343444E410508A5DD1AADD8BD4343524F040853DD",
    INIT_36 => x"08D4DE36ADD8BD554853500408F9DD35ADD8BD534C55500408BCDE34ADD8BD53",
    INIT_37 => x"20DFD9BD415242030869DD3CADD8BD494157430408EDDD37ADD8BD554C555004",
    INIT_38 => x"BD4948420308F8DE219FD9BD4E5242030805DD178DDFD9BD5253420308E0DE16",
    INIT_39 => x"4F4C42030871DE249FD9BD534842030826DF239FD9BD534C42030841DE229FD9",
    INIT_3a => x"4E420308D8DB259FD9BD534342030847DF249FD9BD434342030831DF259FD9BD",
    INIT_3b => x"42030873DF289FD9BD435642030852DF279FD9BD51454203081BDF269FD9BD45",
    INIT_3c => x"03085DDF2B9FD9BD494D42030868DF2A9FD9BD4C50420308C8DE299FD9BD5356",
    INIT_3d => x"089FDF2E9FD9BD5447420308AADF2D9FD9BD544C42030889DF2C9FD9BD454742",
    INIT_3e => x"ECDE243DC1BD3F3C550308CBDF233DC1BD3F3E55030889DE2F9FD9BD454C4203",
    INIT_3f => x"10DF283DC1BD3F53560308C0DF263DC1BD3F3D0208D5DD243DC1BD3F53430308"
    )

    port map (
	  do   => rdata_3,
	  dop(0) => dp(3),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => wdata,
	  dip(0) => dp(3),
	  en   => ce(3),
	  ssr  => rst,
	  we   => we
	);

  RAM4 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0816E02F3DC1BD3F3E02087EDF2C3DC1BD3F3C020804DF2A3DC1BD3F3C300308",
    INIT_01 => x"DD013DC1BD58010894DF003DC1BD44010820E07EC050C901BCC2FFC0BD4F4E02",
    INIT_02 => x"43500208B1DD043DC1BD530108E1DF033DC1BD550108ECDF023DC1BD59010827",
    INIT_03 => x"3DC1BD52434303084BE0093DC1BD42010801E0083DC1BD410108D6DF053DC1BD",
    INIT_04 => x"8118DABD2B2B290308AFDE8018DABD2B29020867E00B3DC1BD5044020839E00A",
    INIT_05 => x"30E08418DABD29010842E08318DABD292D2D030898E08218DABD292D02088EE0",
    INIT_06 => x"0C040CE08B18DABD294402085DE08618DABD2941020879E08518DABD29420208",
    INIT_07 => x"023CDF7EC02029028DD5C3C02820028DD5FFC0BD455A49534548544E45524150",
    INIT_08 => x"12E198C2E6C7B9C902D24EC8E6C76ED6AFC06ED67BCFECE054D4FFC0BD532E02",
    INIT_09 => x"F3D14EC8E6C76ED6AFC06ED67BCFECE054D4FFC0BD532E550306B8E07EC0DBC7",
    INIT_0a => x"7BC20EC9F2C7FDBCC2FFC0BD47534D2E040600E17EC0DBC73AE198C2E6C7B9C9",
    INIT_0b => x"7BC295C6E6C795C626CC7AE16EC2B6C37EC0B0CFB4C60BC47BCFAFC0AEC970E1",
    INIT_0c => x"73654D0A8DD5ECE0AFC0C9C7B0CFB4C626CC26CC76E17BC2D4C895C654C78CE1",
    INIT_0d => x"BCC28DC454D472D4FFC0BD4B4F2E0304F6DF7EC03CD200BCC220232065676173",
    INIT_0e => x"CF4B4F20038DD5DFE16EC26B6F20038DD5D9E17BC295C6DAC4DFE17BC237C901",
    INIT_0f => x"C42BE1FFE17BC237C904BCC28DC4FFE16EC203E1F2E17BC237C902BCC28DC459",
    INIT_10 => x"3CD200BCC264D2E6C795C6CCC492C0D4C895C6CCC40ABCC2AFC037C908BCC28D",
    INIT_11 => x"C53B00CBC2E6C766C5FFC0BD59524555510502A3E07EC02029028DD52CC6CCC4",
    INIT_12 => x"C5FFC0BD4C4C49464552060270E07EC07BCF2CC6BFC400BCC23900CBC281D0A7",
    INIT_13 => x"C0BD3E44524F57050627E17EC0CCC57EC0BFC534E2B5E171E27BC2D4C84EC466",
    INIT_14 => x"07D3F0BCC2A0E298C25CE2D1C6DBC77EC042C891E27BC289C6E6C7D9D3E6C7FF",
    INIT_15 => x"CB580FC401E85886E858891F84A6011F4441455248540604B1E181E26EC2DDC6",
    INIT_16 => x"54C75DC820BCC2AEC989C6E6C7FFC0BD454D414E444E4946080484E0B16E1D03",
    INIT_17 => x"42C8EAE298C26ACB75C7E6C7FEE27BC2E6C795C696CCECE26EC2B0E2F2C74AD3",
    INIT_18 => x"C200C8CCC563E37BC2E6C7EAC6FFC0BD44524F57444E49460804D5E07EC042C8",
    INIT_19 => x"E37BC2D1C6E0C9F2C7DDC642C80ACC76CD42C875C718C795C650CC96CC29E36E",
    INIT_1a => x"C813CDE6C742C863E37BC2E6C7DBC723E398C237C90BC765CDE6C7E6C742C845",
    INIT_1b => x"F2C75BC5F0C3AFC0E6C7D0E2E6C7FFC0BD444E4946040207E37EC039C752CD00",
    INIT_1c => x"A7C4D1C6FFC0BD5453494C44524F572D4843524145530F022EE27EC010E3E0C9",
    INIT_1d => x"C0E6C710E301BCC21DC610C813CDA7C4C3E37BC2F2C7DDC6D0E2E6C7A7C4C2D3",
    INIT_1e => x"7EC03500CBC2A7C4FFC0BD4E4F495443455321080465DE7EC042C8DBC7CCC592",
    INIT_1f => x"E8CCAFC2E6D404E47BC289CD80BCC28000AFC2E6C7FFC0BD2C54494C0404A9E2",
    INIT_20 => x"95C6DAC4FFC0BD4C41524554494C0703C1E07EC0D5E3FDCCBCC2E6D47EC0D5E3",
    INIT_21 => x"E3E8E300C8AFC095C6DAC4FFC0BD4C41524554494C320803DFE07EC0E8E3AFC0",
    INIT_22 => x"FFC0BD3E544947494406064FE17EC04500CBC2FFC0BD4B4F3E0306E3E37EC0E8",
    INIT_23 => x"C296E47BC20EC9F2C710BCC284E47BC20EC9F2C709BCC2E0C930BCC20BC7D1C6",
    INIT_24 => x"B5DF7EC0CCC5DDC6DBC77EC02BC7BFC596E47BC20EC995C6CCC4E6C7E0C907BC",
    INIT_25 => x"CCC488C7D1C6D3E47BC25DE489C6F2C7AFC0E6C7FFC0BD5245424D554E3E0702",
    INIT_26 => x"53554E494D0B0478E27EC0DBC7ACE46EC2B7D201BCC288C7C5CADDC6B2D095C6",
    INIT_27 => x"D201BCC205E57BC2D4C82DBCC289C6F2C705E57BC2E6C7FFC0BD3F4E4749532D",
    INIT_28 => x"88C7E6C7CCC5FFC0BD5245424D554E544F443E0A0455E27EC0CCC57EC0BFC5B7",
    INIT_29 => x"00CBC2E6C7A9E4AEC992C046CE43C9D4C82EBCC289C6F2C733E598C2E6C7B9C9",
    INIT_2a => x"E47EC0A9E4B7D201BCC24700CBC2E6C792C0E2C82EBCC289C6F2C7AFC0E6C747",
    INIT_2b => x"7EC02BC7CCC580E57BC242C817E5D1C6E6E4FFC0BD3F5245424D554E44080629",
    INIT_2c => x"C995C6DAC4AFE57BC2C9C76FE3FFC0BD4C4156450404CCE37EC0BFC586CADDC6",
    INIT_2d => x"E57BC29AC4CBE57BC26BE5A1C6B3C4DBC77EC070C07EC0E8CCABE57BC29EC837",
    INIT_2e => x"71C5FFC0BD504F4F4C2D4B4F0704ADE007D3C3BCC27EC019E4DBC77EC032E4C5",
    INIT_2f => x"D4F8C5FFC0BD544955510402A3DEE8E56EC290E57EE2D6C52CC650CC50CC7CC5",
    INIT_30 => x"CF54E17BCFB0CFA1C6B3C41DE698C260C9E6C7A0D659CFF2D2DBE5AFC234E2F4",
    INIT_31 => x"0526C8FF8310B16E0635042600008310574F52485405026AE3FFE56EC2E5C57B",
    INIT_32 => x"3B00CBC23900CBC2FFC0BD544552505245544E49090496DE07D37EFAE57E0635",
    INIT_33 => x"02DAE47EC0DBC76BE698C289C6E6C7D9D3D6C590E56DE66EC22CC6BFC400BCC2",
    INIT_34 => x"BFC4DDC6F2D255E6AFC2D1C695C6BFC4EAC6A3D2FFC0BD455441554C41564508",
    INIT_35 => x"C292C0FFC0BD444E554F463F060480E67EC030E63B00CBC23900CBC2FBC62CC6",
    INIT_36 => x"C0BD52414843040289E37EC0BAE66FE37EE2D6C5FFC0BD2701028BE507D3F3BC",
    INIT_37 => x"CBE07EC019E4DEE6FFC0BD5D524148435B0603F5E57EC089C6AEC97EE2D6C5FF",
    INIT_38 => x"D429BCC2FFC0BD280103C7E27EC019E437C91FBCC2DEE6FFC0BD4C5254430407",
    INIT_39 => x"29BCC289C6B9C9D7C9A3D244E77BC295C6BFC492C00EC943C495C6BFC446C71F",
    INIT_3a => x"060254E07EC02CC6BFC443C4FFC0BD5C010356E47EC01CE798C25CE292C0D4C8",
    INIT_3b => x"26CC80E77BC20BC703BCC2A7C4D1C6E6C7D0E27EE2D6C5FFC0BD455441455243",
    INIT_3c => x"65520B8DD559CFB7E77BC2DDC600BCC22CC6C0CBAEC989C6F2C7A7C4E6C7DACC",
    INIT_3d => x"C7A7C41DC6B9C9A7C443C98000AFC27BCFB0CFB4C6A7C420676E696E69666564",
    INIT_3e => x"C989C6F2C789C65BC5B9C9A7C42CC600C8A7C42CC696CCA7C495C6E6C7B0E2E6",
    INIT_3f => x"4304045FE77EC0D5E311C16ADBCCC5DACCAEC989C62900CBC2A7C41DC600C843"
    )

    port map (
	  do   => rdata_4,
	  dop(0) => dp(4),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => wdata,
	  dip(0) => dp(4),
	  en   => ce(4),
	  ssr  => rst,
	  we   => we
	);

  RAM5 : RAMB16_S9
    generic map ( 
    INIT_00 => x"D4C3FFC0BD45535255434552070346E46DE76EC2A7C4C2D3A7C4FFC0BD414552",
    INIT_01 => x"C600C843C98000AFC289C6E6C7D4C3FFC0BD4544494804060CE57EC0C8D413CD",
    INIT_02 => x"C01DC600C837C97FBCC289C6E6C7D4C3FFC0BD4C4145564552060629E87EC01D",
    INIT_03 => x"00C843C989C6F2C701BCC2B9C9D4C3FFC0BD4554414944454D4D490902D9E67E",
    INIT_04 => x"454C49504D4F435B09034BE67EC019E4C9E6FFC0BD5D275B0303C7E67EC01DC6",
    INIT_05 => x"C76FE37EE2D6C5FFC0BD454E4F5054534F50080362E57EC0C8D4C9E6FFC0BD5D",
    INIT_06 => x"4F54530506EEE67EC0C8D43500DCC2B3C5D5E3E6D4E6D4D5E87BC29EC8BAE6E6",
    INIT_07 => x"1BBCC20CC2DBC7FDE87BC2D4C8F2C7D6C50CC2DBC7AFC0E6C7F7C1FFC0BD3F50",
    INIT_08 => x"E804D5FCC066E7FFC0BD3A0102ADE87EC0E2C8D6C530E637C9E4BCC2D4C8F2C7",
    INIT_09 => x"DB42CCFCC0AFC2A7C4FFC0BD454D414E4F4E3A070217E77EC0BFCDCCC5BFC52E",
    INIT_0a => x"E6C766E7FFC0BD544E4154534E4F43080201E77EC0D5E3BFCDCCC5CCC504D56A",
    INIT_0b => x"52415608022CE97EC0FDCC3AC17EC0E8CC4FC173E97BC289CD80BCC28000AFC2",
    INIT_0c => x"66E7FFC0BD45554C4156050211E47EC0DACCB3C525C166E7FFC0BD454C424149",
    INIT_0d => x"97E87EC0B4C6AEC9D5C0BDEEC0BD474E495254534F44080414E97EC0E8CC63C1",
    INIT_0e => x"CCC5FDCCE6C76DC801BCC237C9FF00AFC2B2E966E7FFC0BD474E495254530606",
    INIT_0f => x"DDC67EC889C6D1C6AEC9E6C727C2FFC0BD2928244F54050446E87EC0DACCFDCC",
    INIT_10 => x"C989C60BC789C6D1C6AEC9E6C727C2FFC0BD2928244F542B0604FEE77EC0C2D3",
    INIT_11 => x"29282452434E49070464E87EC0A2D363C6DDC6E6C700C8D7C9B4C60BC77EC8E0",
    INIT_12 => x"C21DC6D7C9B4C60BC768EA7BC21BC989C60BC789C6D1C6AEC9E6C727C2FFC0BD",
    INIT_13 => x"DCC2CBC263C170EA40EA0EEAEFE9B2E900007EC02BC7DBC77EC063C6DDC601BC",
    INIT_14 => x"03047CE97EC02700CBC2A7C4E8CCC5C3FFC0BD5453494C584650070413E8F0C2",
    INIT_15 => x"42C8D0EA7BC2D4C895C654C7C5C36CCC95C650CCE6C742CCC9E6FFC0BD584650",
    INIT_16 => x"E907D3E0BCC2B4EA98C2E6C795C650CC7EC0E8CCE8CC42D595C6D7C91FC826CC",
    INIT_17 => x"7EC0A3EA02BCC2FFC0BD4F542B0307DCE87EC0A3EA00BCC2FFC0BD4F540203E9",
    INIT_18 => x"BD53454C424149524156090685EA7EC0A3EA04BCC2FFC0BD52434E49040787E8",
    INIT_19 => x"A7C4C3C6DDC6ACD4FFC0BD455355463C0504E2EA7EC0A2C1DACC7ACC66E7FFC0",
    INIT_1a => x"C2E8CCC3C626CCDACCFEBCC263EB7BC237C90EC9B9C9A7C428C4D4C895C650CC",
    INIT_1b => x"C092C0ABC835EBFFC0BD544958453F0507D3E57EC0D1C626CCE8CCC3C669EB6E",
    INIT_1c => x"C0BFCD01BCC2E8CCE6C7A7C498C27BC2ABC835EBFFC0BD4649020303EB7EC0AF",
    INIT_1d => x"C0BD454C4948570503F2EA94EB6EC26EC2E6D4FFC0BD4441454841050386EB7E",
    INIT_1e => x"A7C495D401BCC2D3CDACD4FFC0BD4E454854040395E97EC012CE01BCC289EBFF",
    INIT_1f => x"C0D5E3BFCD02BCC2A7C4ACD4FFC0BD4E494745420503A9E97EC0D5E32CC600C8",
    INIT_20 => x"7EC0E8CC98C27BC2ABC835EB95D402BCC2D3CDFFC0BD4C49544E550503B8EB7E",
    INIT_21 => x"450403B3E67EC0E8CC6EC2E6D495D402BCC2D3CDFFC0BD4E49414741050304EC",
    INIT_22 => x"29ECFFC0BD54414550455206032FEB7EC0D2EB12CE01BCC2AAEBFFC0BD45534C",
    INIT_23 => x"A4EB7EC0BFCD03BCC2E8CCE6C7A7C407C3E6D4FFC0BD4F44020354EC7EC0D2EB",
    INIT_24 => x"03BCC2D3CDFFC0BD504F4F4C04039FEA71EC6EC225C3E6D4FFC0BD4F443F0303",
    INIT_25 => x"FFC0BD504F4F4C2B05033EEC7EC02CC600C8A7C4E8CC26CCE6C73DC3E6D495D4",
    INIT_26 => x"EC7BC295D4CCC5D3CDFFC0BD3B010323ECA6EC6EC262C3E6D495D403BCC2D3CD",
    INIT_27 => x"5202074FE77EC0D2EB7EC0E6D4FFC0BD7D010770EB7EC0F4D47EC0E6D44DE8E3",
    INIT_28 => x"ABC835EBFFC0BD45523F0307D2EC7EC0E8CC42CC13CDD4C36EC2E6D4FFC0BD45",
    INIT_29 => x"4E4F4F4406042AE67EC0D2EB01EDFFC0BD7D4552030715EB08ED6EC27BC298C2",
    INIT_2a => x"A1E47EC01DC62D00CBC2E6C7B9C91DC654C7B9C95BC589C6D5C0BDEEC0BD594C",
    INIT_2b => x"45EDBD594C4E4F040281EC7EC01DC6F0C389C6D5C0BDEEC0BD434F564F440504",
    INIT_2c => x"046AEDBD454449534E49060050E980ED026AEDBD4854524F46050067EC000000",
    INIT_2d => x"EDBD52454C424D45535341090007EA9FED066AEDBD41525458450500EEEC8FED",
    INIT_2e => x"D7C902BCC289C6E6C7A7C3A7C4FFC0BD5453494C44524F570802B7ECAEED086A",
    INIT_2f => x"C80EC9F0C34CC5FFC0BD4F534C410400C7ED7EC089C62300CBC2E6C7E8CCFDCC",
    INIT_30 => x"455250080061ED7EC01DC6F0C32D00DCC2FFBCC289C6F0C330E637C9CFBCC2AB",
    INIT_31 => x"ED7EC02D00F0C230E637C9CEBCC2ABC80EC95BC5AEC9F0C3FFC0BD53554F4956",
    INIT_32 => x"470B00A5ED7EC01DC65BC589C6F0C3FFC0BD534E4F4954494E494645440B003B",
    INIT_33 => x"45525255432D5445530B0038EA7EC089C65BC5FFC0BD544E45525255432D5445",
    INIT_34 => x"C889C654C7A7C3FFC0BD454D414E434F560704FEEC7EC01DC65BC5FFC0BD544E",
    INIT_35 => x"46C79BEE98C2E6C795C6AEC97EC037C91FBCC2B4C628CD6CCC42C8B4EE7BC2D4",
    INIT_36 => x"524544524F0500F1ED7EC0B0CF96EEFFC0BD434F562E0406CDEB7EC03F017DD5",
    INIT_37 => x"8DD5F4EE3DC37BCFCEEEB4C6FEEE07C300BCC2E0C9F2C75BC5F0C3ECE0FFC0BD",
    INIT_38 => x"C0F6ED8CEDF6EDABED7DEDFFC0BD4853455246050086ED7EC0CEEE89C6203A02",
    INIT_39 => x"0704DAEE7EC067EDDBC7D0ED66E7FFC0BD5952414C554241434F560A0693EC7E",
    INIT_3a => x"8FC8E0C93AC595C688C366EF07C303BCC223BCC2CCC5FFC0BD41464E504F5421",
    INIT_3b => x"D1C6FFC0BD4C494154525543070476EE7EC02900CBC2D7C93AC556EF62C3B3C5",
    INIT_3c => x"524F4628070424EF7EC02BC784EF98C289CD75C7E6C795C6D7C90BC78AEF6EC2",
    INIT_3d => x"C52CC688C37BEFFDBCC295C688C3C5EF07C303BCC223BCC2A7C4FFC0BD544547",
    INIT_3e => x"FEBCC2C5C32500CBC27BEF02BCC2B6C32300CBC27BEF01BCC2A7C3B2EF62C3B3",
    INIT_3f => x"C67EE2D6C5FFC0BD544547524F4606021CEE7EC047EFDACCE0C92700CBC27BEF"
    )

    port map (
	  do   => rdata_5,
	  dop(0) => dp(5),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => wdata,
	  dip(0) => dp(5),
	  en   => ce(5),
	  ssr  => rst,
	  we   => we
	);

  RAM6 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0EC9F2C7A7C4E0C937C902BCC265CD00C896CCE6C728CDBAE699E389C65BC5B4",
    INIT_01 => x"8000AFC289C6D4C3FFC0BD45564F4D455206068EEE7EC0A3EF30E637C9F1BCC2",
    INIT_02 => x"52454B52414D4F4408042EF00BF06EC27BCFB0CFB4C6E6C7D4C34DE8AFC037C9",
    INIT_03 => x"A2D3AEC9E0C9F2C75BC52D00CBC2E6C7B4C626CCA3EF95C6E6C7D5C0BDEEC0BD",
    INIT_04 => x"C5A7C4FDCCE6C7F0C3E8CC60F066E7A7C4FFC0BD52454B52414D0602B4ED7EC0",
    INIT_05 => x"D1C695C6BFC4FFC0BD57454E4104063FEF7EC0A2D3DACCE6C7AEC9E0C9F0C35B",
    INIT_06 => x"C9E6C7F5F07BC2C9C737C9F2C86FE330E637C9E0BCC2ABC889C6E6C7D9D3D6C5",
    INIT_07 => x"EE7EC08CF02CC6BFC4DDC670C0F5F07BC2C9C737C9D4C860F0AFC26CCC95C6AE",
    INIT_08 => x"95C682C44300DCC20008AFC24300CBC200F8AFC2FFC0BD4D454D49482106045E",
    INIT_09 => x"0602C1E97EC014F17BC2E2C860C92CC682C4F2C795C682C42CC682C460C9E6C7",
    INIT_0a => x"1F4F444C4F43040695ED7EC0E0C9A7C4E0C920BCC282C4FFC0BD444553554E55",
    INIT_0b => x"CBC200BCC247EF09F19ACB65BCC200BCC23AC5FFC0BDFE01CE06357E01CE108B",
    INIT_0c => x"7279706F431F8DD559CF54E100BCC259CFE4C17FBCC24EEE12EFDBC71DD52F00",
    INIT_0d => x"531D8DD559CF67672D6874726F46204343482035303032202963282074686769",
    INIT_0e => x"82C459CF72656E6265754820736E61482079622074726F702039306D65747379",
    INIT_0f => x"442806049BEFFAE559CF59CF4D415220426B20078DD53CD209BCC288C90ABCC2",
    INIT_10 => x"D4F2C7CCC5D3CDFFC0BD3E53454F440503FDF17EC03DCDDDC6FFC0BD3E53454F",
    INIT_11 => x"BCC266E7FFC0BD45444F43040215ED7EC0D5E36ADBD5C0AFC204F2E6D4BFCD95",
    INIT_12 => x"CCC5D3CDFFC0BD45444F433B05033FF17EC0BFCD05BCC2BFC52EE8BEEDDACCFD",
    INIT_13 => x"C016E9FFC0BD3A52454F4405062BED7EC0F4D4BEED04F2E6D4BFCD05BCC295D4",
    INIT_14 => x"C0DACC03BCC239F2FFC0BD45444F4352454F44080642EE7EC06ADBD5C0AFC2EB",
    INIT_15 => x"EE4DE8BFF27BC295D405BCC2D3CDFFC0BD45444F432D444E450808B2F07EC0EB",
    INIT_16 => x"414E45060673EF7EC02CC6AEC9FFC0BD524F5443455621070634F27EC0F6ED25",
    INIT_17 => x"3BBCC2FFC0BD454C424153494407060CEF7EC01DC600C87EBCC2FFC0BD454C42",
    INIT_18 => x"EF7EC02CC6BFC437C9E2E895C6BFC4FFC0BD594E414D0406A6F27EC01DC600C8",
    INIT_19 => x"43C9E2E8D4C80BC73700CBC200BCC2D1C6AEC937C4FFC0BD53454D49540506F1",
    INIT_1a => x"5344524F570B0409F37EC02CC6BFC400BCC23700CBC2DDC67EC02BC748F37BC2",
    INIT_1b => x"C2D4C876CD54C783F37BC2E6C795C696CC71F36EC200C8FFC0BD52455050494B",
    INIT_1c => x"C7D7C924BCC25CC43CC61DD5FFC0BD5344524F5728060422F37EC042C86FF37B",
    INIT_1d => x"88C370C0A1C65CC488C3C8F307C354C79ACB20BCC2F2C703BCC2E0C920BCC2E6",
    INIT_1e => x"7BC295C688C304F407C375C7FFBCC2CCC5D1C600BCC259CFB6F362C3B3C52CC6",
    INIT_1f => x"B3C588C3E0C93AC595C688C346C7FEF37BC20EC9E0C93AC595C688C3F2C7FEF3",
    INIT_20 => x"C03CD200BCC2ECE0DDC659CF46C7DBC721F47BC243C9E2E846CE42C8DAF362C3",
    INIT_21 => x"BCC2E6C7B4C6E6C795C6E6C7D1C6AEC9DDC659CF2EF47BC20EC968C43CBCC27E",
    INIT_22 => x"C65CC496CC7BCFB0CF48CF7EBCC237C91FBCC255F46EC2D6C54DF47BC228C920",
    INIT_23 => x"F366F3AFC289C6F0C3FFC0BD5344524F57050053F2CFF36EC22CC600C870C0A1",
    INIT_24 => x"EBEB7EC091F370C0AFC295C6AFC2FFC0BD5344524F574C4C410806DCF27EC091",
    INIT_25 => x"44412E0404A1F47EC01DC65CC442C873D146CEFF00AFC2FFC0BD21522E580404",
    INIT_26 => x"3CD289C65CC4FFC0BD455459422E050457F07EC026D2C4C989C65CC4FFC0BD52",
    INIT_27 => x"74F27EC048CF6DC8D6C537C928C97FBCC2E6C7FFC0BD4353412E0404C9EE7EC0",
    INIT_28 => x"C921F57BC228C906BCC2E6C75DC810BCC295C6CCC4A6F4FFC0BD504D55440402",
    INIT_29 => x"D7C988C3E6C74AF507C300BCC20BC77BCFC1F459CFE6C700C8D7C9F2C7D1C6C4",
    INIT_2a => x"D557F53DC3EAF4B4C65FF507C300BCC20BC77C018DD53AF53DC37BCFD7F489C6",
    INIT_2b => x"0504C8F27EC02BC746C729F57BC243C9E2E80EC90BC7E0C900C854C7207C028D",
    INIT_2c => x"E6C7B9C900C837C989CDA7C43AC5F2C70EC9F2C70003AFC2FFC0BD3F3F414643",
    INIT_2d => x"C789C6F2C7DDC6B9C9D1C601BCC2AFC0E6C737C937C989CD7FBCC221BCC289C6",
    INIT_2e => x"C9F2C7D6C5AEC9E5F57BC289CD7FBCC221BCC27EC0F2C846C7CDF57BC2D4C854",
    INIT_2f => x"AFC0E6C737C985F5E6C7FFC0BD3F414643040478ED7EC0CCC546C7B5F57BC237",
    INIT_30 => x"B9C922F698C2E6C795C696CCAFC0E6C737C9ABC828C976CDF2C789C6A7C328CD",
    INIT_31 => x"F2F27EC0CCC5DBC77EC085F513CD38F67BC289CD20BCC200BCC289C6E6C77EC0",
    INIT_32 => x"CFB4C628CDB0CF18C7EAC620202D2D2020067DD5E6C7FFC0BD444145482E0504",
    INIT_33 => x"CD2072656F64058DD5E6C785F67BC2F3F5E6C76CCC95C6AEC9E6C7B0CF18C7B0",
    INIT_34 => x"2E0604BCF47EC064726F5720058DD5CEEE76CD28CDB0CFFBC6DBC7B0CFB4C628",
    INIT_35 => x"B0CFB4C628CD8ECFD7C904BCC2C4C9C4C937C901BCC2F2C7FFC0BD4E454B4F54",
    INIT_36 => x"F4E6C7B4C6E6C7203A028DD5C1F4E6C759CFFFC0BD4D4F43454405049EF67EC0",
    INIT_37 => x"01BCC2F2C7D6C5C1F495C6E6C77BCFEAF47BCFD7F4E6C789C67BCFEAF47BCFD7",
    INIT_38 => x"C77EC0AEC947F6E6C71FF77BC2F3F5E6C77BCF48CFD7C90EBCC20BF77BC237C9",
    INIT_39 => x"C992C0F3F595C6E6C792C0F3F5E6C7AEC9A5F695C6E6C743F77BC2F3F595C6E6",
    INIT_3a => x"7EC0DBC754F77BC2E2E8CBF6A6F4FFC0BD4545534D040686F47EC0AEC97EC0AE",
    INIT_3b => x"BDEEC0BD4553414246464F4408048CF27EC04FF7C9E6FFC0BD45455303026EF4",
    INIT_3c => x"30E62CC6CCC4DDC6F2D290E5AFC27EE2D6C52CC6CCC489C6D1C695C6CCC4D5C0",
    INIT_3d => x"BD58480201D1F47EC06EE8FDCC7CF766E7FFC0BD455341424646060401F57EC0",
    INIT_3e => x"4E4548545B06017FF5027FF7BD4E420201C6F70A7FF7BD4D4402018AF3107FF7",
    INIT_3f => x"DBC700F86EC2FFC0BD5D4C414E4F495449444E4F435B0D0463F77EC0FFC0BD5D"
    )

    port map (
	  do   => rdata_6,
	  dop(0) => dp(6),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => wdata,
	  dip(0) => dp(6),
	  en   => ce(6),
	  ssr  => rst,
	  we   => we
	);

  RAM7 : RAMB16_S9
    generic map ( 
    INIT_00 => x"54C74AD354C7B7D201BCC2B4C6FEF77BC2D4C85BBCC289C6AEC9E6C77EE2D6C5",
    INIT_01 => x"5D45534C45057DD554C7FAF76EC2AFC046C736F898C273D35D4E454854057DD5",
    INIT_02 => x"46C768F898C273D35D4649037DD554C7FAF76EC2AFC0C9C746C750F898C273D3",
    INIT_03 => x"F7FAF76EC2AEC9E6C77BF898C273D35D4441454841067DD5FAF76EC2AEC9E6C7",
    INIT_04 => x"C0BD5D44414548415B0701EEF57EC0F7F700BCC2FFC0BD5D45534C455B0601DA",
    INIT_05 => x"C2FFC0BD534D020202F17EC089F892C0FFC0BD5D46495B040185F07EC089F8FF",
    INIT_06 => x"0188A8F813D17EC0C6F83DC3D0F83DC3D4F807C300BCC212BCC2D8F825C300BC",
    INIT_07 => x"B4C6D9D3D6C500BCC2FFC0BD4745520309BCF77EC03300CBC200BCC2FFC0BD23",
    INIT_08 => x"F8E6D4E8E342D5DBC707F93DC3DDC643C9D1C600C8FBD6B4C617F925C300BCC2",
    INIT_09 => x"BD2950440308C5F67EC0E1F8FF00AFC2FFC0BD4745524C4C4106084AF77EC0E1",
    INIT_0a => x"73F77EC0D0D68900AFC200C8FFC0BD2923020882F87EC03300CBC210BCC2FFC0",
    INIT_0b => x"18C4FFC0BD5D5B02084EF97EC08D00AFC23300CBC220BCC2FFC0BD2943500308",
    INIT_0c => x"7EC0D7C910BCC2B8D6D4C88000AFC237C99D00AFC2E6C7A0F97BC2D4C820BCC2",
    INIT_0d => x"C4FDCC00BCC2FDCCFFC0BD4649028896F886EB7EC09F00AFC23300CBC220BCC2",
    INIT_0e => x"F4CDEB7EC0B5F920BCC2FFC0BD44414548410588B2F9A4EB7EC0BFCD06BCC2A7",
    INIT_0f => x"C8B8D6ABC886D6E6C7E0C9F2C7A7C495D406BCC2D3CDFFC0BD4E4548540488E5",
    INIT_10 => x"04EC7EC0BFCD07BCC2A7C4FFC0BD4E4947454205883BF9EBEB7EC01DC6B9C900",
    INIT_11 => x"D6E6C7E0C9AEC9A7C4FDCC00C895D407BCC2D3CDFFC0BD4C49544E55058878F9",
    INIT_12 => x"3EEC7EC029FA20BCC2FFC0BD4E49414741058823FA23EC7EC0FDCCB8D6ABC886",
    INIT_13 => x"45504552068841F654EC7EC0E7F912CE01BCC2D3F9FFC0BD45534C4504885AF3",
    INIT_14 => x"12CE01BCC2B5F9FFC0BD454C49485705884EFAB8EB7EC0E7F954FAFFC0BD5441",
    INIT_15 => x"2D444345530B0690FA7EC0ACDA7BF99CE044E0FFC0BD5458454E0408D0F77EC0",
    INIT_16 => x"484749482D535345524444412D44434553110626F940B152C1BD535554415453",
    INIT_17 => x"530A06B9F800B252C1BD455341422D4D41522D444345530D06CDF941B152C1BD",
    INIT_18 => x"544154532D444345532E0C06E2F97EC002D2A7C4FFC0BD54524154532D444345",
    INIT_19 => x"088DD5B5F9ABC837C901BCC2E6C789C6C6FA203A44434553068DD5FFC0BD5355",
    INIT_1a => x"C903BCC288C901BCC2E7F920444550504F5453088DD568FA20474E494E4E5552",
    INIT_1b => x"D5B5F9D4C801BCC2E6C7E7F9474E494E4E5552078DD5B5F9D4C800BCC2E6C737",
    INIT_1c => x"F9D4C803BCC2E7F94347028DD5B5F9D4C802BCC2E6C7E7F94445544C4148068D",
    INIT_1d => x"BD454741502D444345532E0A0610F27EC059CFE7F94E574F4E4B4E55078DD5B5",
    INIT_1e => x"4553080659F17EC02CC6CCC406F50001AFC2F6FA77D295C6CCC41DC6E0FAFFC0",
    INIT_1f => x"6E61206874726F467369614D0F000000007EC002D2A7C4FFC0BD444E452D4443",
    INIT_20 => x"6B636174530F03FCFCFF776F6C667265766F206B636174530EEFFBFDFF313036",
    INIT_21 => x"6E4F0E2AFCF2FF646E69662074276E61430A16FCF3FF776F6C667265646E7520",
    INIT_22 => x"450C4CFCF0FF6465746365746F72500939FCF1FF676E696C69706D6F6320796C",
    INIT_23 => x"FF726F727265206572757463757274530F5AFCEAFF7475706E6920666F20646E",
    INIT_24 => x"6E2064696C61766E49157FFCE0FF747075727265746E6920726573550E6BFCE4",
    INIT_25 => x"766F20726564726F206863726165531592FCCFFF746E656D7567726120656D61",
    INIT_26 => x"6F6C667265646E7520726564726F2068637261655316ACFCCEFF776F6C667265",
    INIT_27 => x"72207369204553414218E1FCC2FF3F73696874207327746168570CC6FCC3FF77",
    INIT_28 => x"72646461206C6167656C6C4917F2FCC1FF6C616D69636564206F742074657365",
    INIT_29 => x"00000000000000000000000000000000E2C000000065646F6D20676E69737365",
    INIT_2a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3f => x"5EF1640061005E005B005800550000C000000000000000000000000000000000"
    )

    port map (
	  do   => rdata_7,
	  dop(0) => dp(7),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => wdata,
	  dip(0) => dp(7),
	  en   => ce(7),
	  ssr  => rst,
	  we   => we
	);

my_rom_16k : process ( cs, rw, addr,
                       rdata_0, rdata_1, rdata_2, rdata_3,
                       rdata_4, rdata_5, rdata_6, rdata_7)
begin
	 we <= not rw;
	 
	 case addr(13 downto 11) is
	 when "000" =>
	     rdata <= rdata_0;
	 when "001" =>
	     rdata <= rdata_1;
	 when "010" =>
	     rdata <= rdata_2;
	 when "011" =>
	     rdata <= rdata_3;
	 when "100" =>
	     rdata <= rdata_4;
	 when "101" =>
	     rdata <= rdata_5;
	 when "110" =>
	     rdata <= rdata_6;
	 when "111" =>
	     rdata <= rdata_7;
	 when others =>
	     null;
    end case;

    ce(0)  <= cs and not( addr(13) ) and not( addr(12) ) and not( addr(11) );
    ce(1)  <= cs and not( addr(13) ) and not( addr(12) ) and      addr(11)  ;
    ce(2)  <= cs and not( addr(13) ) and      addr(12)   and not( addr(11) );
    ce(3)  <= cs and not( addr(13) ) and      addr(12)   and      addr(11)  ;
    ce(4)  <= cs and      addr(13)   and not( addr(12) ) and not( addr(11) );
    ce(5)  <= cs and      addr(13)   and not( addr(12) ) and      addr(11)  ;
    ce(6)  <= cs and      addr(13)   and      addr(12)   and not( addr(11) );
    ce(7)  <= cs and      addr(13)   and      addr(12)   and      addr(11)  ;

end process;

end architecture rtl;

